module instmem_aes128_m1 (a,inst);
    input  [31:0] a;
    output [31:0] inst;
    wire   [31:0] rom [0:511];
    // aes_128_enc_key_schedule:
    assign rom[9'h000] = 32'b00000100100000000000001010010011; // la  t0,  initial_key
    assign rom[9'h001] = 32'b00000000000000101010010110000011; // lw  a1,   0(t0) 
    assign rom[9'h002] = 32'b00000000010000101010011000000011; // lw  a2,   4(t0) 
    assign rom[9'h003] = 32'b00000000100000101010011010000011; // lw  a3,   8(t0) 
    assign rom[9'h004] = 32'b00000000110000101010011100000011; // lw  a4,  12(t0) 
    assign rom[9'h005] = 32'b00000101100000000000010100010011; // la    a0,  round_key
    assign rom[9'h006] = 32'b00001010000001010000001010010011; // addi  t0,  a0,  160
    assign rom[9'h007] = 32'b00000000000000000000001100010011; // la    t1,  aes_round_const
    // aes_128_enc_ks_l0:
    assign rom[9'h008] = 32'b00000000101101010010000000100011; // sw  a1,   0(a0)
    assign rom[9'h009] = 32'b00000000110001010010001000100011; // sw  a2,   4(a0) 
    assign rom[9'h00a] = 32'b00000000110101010010010000100011; // sw  a3,   8(a0)
    assign rom[9'h00b] = 32'b00000000111001010010011000100011; // sw  a4,  12(a0)
    assign rom[9'h00c] = 32'b00000010010101010000110001100011; // beq  a0,  t0,  aes_128_enc_ks_finish
    assign rom[9'h00d] = 32'b00000001000001010000010100010011; // addi  a0,  a0,  16
    assign rom[9'h00e] = 32'b00000000000000110100001110000011; // lbu   t2,  0(t1)
    assign rom[9'h00f] = 32'b00000000010000110000001100010011; // addi  t1,  t1,  4
    assign rom[9'h010] = 32'b00000000011101011100010110110011; // xor   a1,  a1,  t2
    assign rom[9'h011] = 32'b00000001100001110001010000010011; // slli  s0,  a4,  24
    assign rom[9'h012] = 32'b00000000100001110101010010010011; // srli  s1,  a4,  8
    assign rom[9'h013] = 32'b00000000100101000110010000110011; // or    s0,  s0,  s1   
    assign rom[9'h014] = 32'b00000010000001000000010001111111; // subbytes  s0,  s0
    assign rom[9'h015] = 32'b00000000100001011100010110110011; // xor  a1,  a1,  s0
    assign rom[9'h016] = 32'b00000000101101100100011000110011; // xor  a2,  a2,  a1
    assign rom[9'h017] = 32'b00000000110001101100011010110011; // xor  a3,  a3,  a2
    assign rom[9'h018] = 32'b00000000110101110100011100110011; // xor  a4,  a4,  a3
    assign rom[9'h019] = 32'b11111011110111111111000001101111; // j   aes_128_enc_ks_l0
    // aes_128_enc_ks_finish:
    assign rom[9'h01a] = 32'b00000101100000000000010100010011; // la  a0,  round_key
    // aes_128_encrypt:
    assign rom[9'h01b] = 32'b00000000101000000000011110010011; // li    a5,  10
    assign rom[9'h01c] = 32'b00000000010001111001100000010011; // slli  a6,  a5,  4
    assign rom[9'h01d] = 32'b00000000101010000000100000110011; // add   a6,  a6,  a0
    assign rom[9'h01e] = 32'b00000010100000000000100010010011; // la    a7,  input_block
    assign rom[9'h01f] = 32'b00000000000010001010100100000011; // lw    s2,   0(a7)
    assign rom[9'h020] = 32'b00000000010010001010100110000011; // lw    s3,   4(a7)
    assign rom[9'h021] = 32'b00000000100010001010101000000011; // lw    s4,   8(a7)
    assign rom[9'h022] = 32'b00000000110010001010101010000011; // lw    s5,  12(a7)
    assign rom[9'h023] = 32'b00000000000001010010101100000011; // lw    s6,  0(a0)
    assign rom[9'h024] = 32'b00000000010001010010101110000011; // lw    s7,  4(a0)
    assign rom[9'h025] = 32'b00000000100001010010110000000011; // lw    s8,  8(a0)
    assign rom[9'h026] = 32'b00000000110001010010110010000011; // lw    s9, 12(a0)
    assign rom[9'h027] = 32'b00000001011010010100100100110011; // xor   s2,  s2,  s6
    assign rom[9'h028] = 32'b00000001011110011100100110110011; // xor   s3,  s3,  s7
    assign rom[9'h029] = 32'b00000001100010100100101000110011; // xor   s4,  s4,  s8
    assign rom[9'h02a] = 32'b00000001100110101100101010110011; // xor   s5,  s5,  s9
    assign rom[9'h02b] = 32'b00000001000001010000010100010011; // addi  a0,  a0,  16
    assign rom[9'h02c] = 32'b00001111111100000000000110010011; // li    gp,  0xFF
    // aes_enc_block_loop:
    assign rom[9'h02d] = 32'b00000010000010010000101101111111; // subbytes  s6,  s2
    assign rom[9'h02e] = 32'b00000010000010011000101111111111; // subbytes  s7,  s3
    assign rom[9'h02f] = 32'b00000010000010100000110001111111; // subbytes  s8,  s4
    assign rom[9'h030] = 32'b00000010000010101000110011111111; // subbytes  s9,  s5
    assign rom[9'h031] = 32'b00000000001110110111100100110011; // and   s2,   s6,   gp
    assign rom[9'h032] = 32'b00000000001110111111100110110011; // and   s3,   s7,   gp
    assign rom[9'h033] = 32'b00000000001111000111101000110011; // and   s4,   s8,   gp
    assign rom[9'h034] = 32'b00000000001111001111101010110011; // and   s5,   s9,   gp
    assign rom[9'h035] = 32'b00000000100000011001110100010011; // slli  s10,  gp,   0x8
    assign rom[9'h036] = 32'b00000001101010111111110110110011; // and   s11,  s7,   s10
    assign rom[9'h037] = 32'b00000001101110010110100100110011; // or    s2,   s2,   s11
    assign rom[9'h038] = 32'b00000001101011000111110110110011; // and   s11,  s8,   s10
    assign rom[9'h039] = 32'b00000001101110011110100110110011; // or    s3,   s3,   s11
    assign rom[9'h03a] = 32'b00000001101011001111110110110011; // and   s11,  s9,   s10
    assign rom[9'h03b] = 32'b00000001101110100110101000110011; // or    s4,   s4,   s11
    assign rom[9'h03c] = 32'b00000001101010110111110110110011; // and   s11,  s6,   s10
    assign rom[9'h03d] = 32'b00000001101110101110101010110011; // or    s5,   s5,   s11
    assign rom[9'h03e] = 32'b00000000100011010001110100010011; // slli  s10,  s10,  0x8
    assign rom[9'h03f] = 32'b00000001101011000111110110110011; // and   s11,  s8,   s10
    assign rom[9'h040] = 32'b00000001101110010110100100110011; // or    s2,   s2,   s11
    assign rom[9'h041] = 32'b00000001101011001111110110110011; // and   s11,  s9,   s10
    assign rom[9'h042] = 32'b00000001101110011110100110110011; // or    s3,   s3,   s11
    assign rom[9'h043] = 32'b00000001101010110111110110110011; // and   s11,  s6,   s10
    assign rom[9'h044] = 32'b00000001101110100110101000110011; // or    s4,   s4,   s11
    assign rom[9'h045] = 32'b00000001101010111111110110110011; // and   s11,  s7,   s10
    assign rom[9'h046] = 32'b00000001101110101110101010110011; // or    s5,   s5,   s11
    assign rom[9'h047] = 32'b00000000100011010001110100010011; // slli  s10,  s10,  0x8
    assign rom[9'h048] = 32'b00000001101011001111110110110011; // and   s11,  s9,   s10
    assign rom[9'h049] = 32'b00000001101110010110100100110011; // or    s2,   s2,   s11
    assign rom[9'h04a] = 32'b00000001101010110111110110110011; // and   s11,  s6,   s10
    assign rom[9'h04b] = 32'b00000001101110011110100110110011; // or    s3,   s3,   s11
    assign rom[9'h04c] = 32'b00000001101010111111110110110011; // and   s11,  s7,   s10
    assign rom[9'h04d] = 32'b00000001101110100110101000110011; // or    s4,   s4,   s11
    assign rom[9'h04e] = 32'b00000001101011000111110110110011; // and   s11,  s8,   s10
    assign rom[9'h04f] = 32'b00000001101110101110101010110011; // or    s5,   s5,   s11
    assign rom[9'h050] = 32'b00000100000010010000100101111111; // mixColumns  s2,  s2
    assign rom[9'h051] = 32'b00000100000010011000100111111111; // mixColumns  s3,  s3
    assign rom[9'h052] = 32'b00000100000010100000101001111111; // mixColumns  s4,  s4
    assign rom[9'h053] = 32'b00000100000010101000101011111111; // mixColumns  s5,  s5
    assign rom[9'h054] = 32'b00000000000001010010101100000011; // lw    s6,   0(a0)
    assign rom[9'h055] = 32'b00000000010001010010101110000011; // lw    s7,   4(a0)
    assign rom[9'h056] = 32'b00000000100001010010110000000011; // lw    s8,   8(a0)
    assign rom[9'h057] = 32'b00000000110001010010110010000011; // lw    s9,  12(a0)
    assign rom[9'h058] = 32'b00000001011010010100100100110011; // xor   s2,  s2,  s6
    assign rom[9'h059] = 32'b00000001011110011100100110110011; // xor   s3,  s3,  s7
    assign rom[9'h05a] = 32'b00000001100010100100101000110011; // xor   s4,  s4,  s8
    assign rom[9'h05b] = 32'b00000001100110101100101010110011; // xor   s5,  s5,  s9
    assign rom[9'h05c] = 32'b00000001000001010000010100010011; // addi  a0,  a0,  16
    assign rom[9'h05d] = 32'b11110101000001010001000011100011; // bne   a0,  a6,  aes_enc_block_loop
    // aes_enc_block_finish:
    assign rom[9'h05e] = 32'b00000010000010010000101101111111; // subbytes  s6,   s2
    assign rom[9'h05f] = 32'b00000010000010011000101111111111; // subbytes  s7,   s3
    assign rom[9'h060] = 32'b00000010000010100000110001111111; // subbytes  s8,   s4
    assign rom[9'h061] = 32'b00000010000010101000110011111111; // subbytes  s9,   s5 
    assign rom[9'h062] = 32'b00000000001110110111100100110011; // and   s2,   s6,   gp
    assign rom[9'h063] = 32'b00000000001110111111100110110011; // and   s3,   s7,   gp
    assign rom[9'h064] = 32'b00000000001111000111101000110011; // and   s4,   s8,   gp
    assign rom[9'h065] = 32'b00000000001111001111101010110011; // and   s5,   s9,   gp
    assign rom[9'h066] = 32'b00000000100000011001110100010011; // slli  s10,  gp,   0x8
    assign rom[9'h067] = 32'b00000001101010111111110110110011; // and   s11,  s7,   s10
    assign rom[9'h068] = 32'b00000001101110010110100100110011; // or    s2,   s2,   s11
    assign rom[9'h069] = 32'b00000001101011000111110110110011; // and   s11,  s8,   s10
    assign rom[9'h06a] = 32'b00000001101110011110100110110011; // or    s3,   s3,   s11
    assign rom[9'h06b] = 32'b00000001101011001111110110110011; // and   s11,  s9,   s10
    assign rom[9'h06c] = 32'b00000001101110100110101000110011; // or    s4,   s4,   s11
    assign rom[9'h06d] = 32'b00000001101010110111110110110011; // and   s11,  s6,   s10
    assign rom[9'h06e] = 32'b00000001101110101110101010110011; // or    s5,   s5,   s11
    assign rom[9'h06f] = 32'b00000000100011010001110100010011; // slli  s10,  s10,  0x8
    assign rom[9'h070] = 32'b00000001101011000111110110110011; // and   s11,  s8,   s10
    assign rom[9'h071] = 32'b00000001101110010110100100110011; // or    s2,   s2,   s11
    assign rom[9'h072] = 32'b00000001101011001111110110110011; // and   s11,  s9,   s10
    assign rom[9'h073] = 32'b00000001101110011110100110110011; // or    s3,   s3,   s11
    assign rom[9'h074] = 32'b00000001101010110111110110110011; // and   s11,  s6,   s10
    assign rom[9'h075] = 32'b00000001101110100110101000110011; // or    s4,   s4,   s11
    assign rom[9'h076] = 32'b00000001101010111111110110110011; // and   s11,  s7,   s10
    assign rom[9'h077] = 32'b00000001101110101110101010110011; // or    s5,   s5,   s11
    assign rom[9'h078] = 32'b00000000100011010001110100010011; // slli  s10,  s10,  0x8
    assign rom[9'h079] = 32'b00000001101011001111110110110011; // and   s11,  s9,   s10
    assign rom[9'h07a] = 32'b00000001101110010110100100110011; // or    s2,   s2,   s11
    assign rom[9'h07b] = 32'b00000001101010110111110110110011; // and   s11,  s6,   s10
    assign rom[9'h07c] = 32'b00000001101110011110100110110011; // or    s3,   s3,   s11
    assign rom[9'h07d] = 32'b00000001101010111111110110110011; // and   s11,  s7,   s10
    assign rom[9'h07e] = 32'b00000001101110100110101000110011; // or    s4,   s4,   s11
    assign rom[9'h07f] = 32'b00000001101011000111110110110011; // and   s11,  s8,   s10
    assign rom[9'h080] = 32'b00000001101110101110101010110011; // or    s5,   s5,   s11
    assign rom[9'h081] = 32'b00000000000001010010101100000011; // lw   s6,   0(a0)
    assign rom[9'h082] = 32'b00000000010001010010101110000011; // lw   s7,   4(a0)
    assign rom[9'h083] = 32'b00000000100001010010110000000011; // lw   s8,   8(a0)
    assign rom[9'h084] = 32'b00000000110001010010110010000011; // lw   s9,  12(a0)
    assign rom[9'h085] = 32'b00000001011010010100100100110011; // xor  s2,  s2,  s6
    assign rom[9'h086] = 32'b00000001011110011100100110110011; // xor  s3,  s3,  s7
    assign rom[9'h087] = 32'b00000001100010100100101000110011; // xor  s4,  s4,  s8
    assign rom[9'h088] = 32'b00000001100110101100101010110011; // xor  s5,  s5,  s9
    assign rom[9'h089] = 32'b00000011100000000000100010010011; // la   a7,  output_block
    assign rom[9'h08a] = 32'b00000001001010001010000000100011; // sw   s2,   0(a7)
    assign rom[9'h08b] = 32'b00000001001110001010001000100011; // sw   s3,   4(a7)
    assign rom[9'h08c] = 32'b00000001010010001010010000100011; // sw   s4,   8(a7)
    assign rom[9'h08d] = 32'b00000001010110001010011000100011; // sw   s5,  12(a7)
    // aes_128_decrypt:
    assign rom[9'h08e] = 32'b00000101100000000000100000010011; // la  a6,  round_key
    assign rom[9'h08f] = 32'b00000000101000000000011110010011; // li    a5,  10
    assign rom[9'h090] = 32'b00000000010001111001010100010011; // slli  a0,  a5,  4
    assign rom[9'h091] = 32'b00000001000001010000010100110011; // add   a0,  a0,  a6
    assign rom[9'h092] = 32'b00000011100000000000100010010011; // la    a7,  output_block
    assign rom[9'h093] = 32'b00000000000010001010100100000011; // lw    s2,   0(a7)
    assign rom[9'h094] = 32'b00000000010010001010100110000011; // lw    s3,   4(a7)
    assign rom[9'h095] = 32'b00000000100010001010101000000011; // lw    s4,   8(a7)
    assign rom[9'h096] = 32'b00000000110010001010101010000011; // lw    s5,  12(a7)
    assign rom[9'h097] = 32'b00000000000001010010101100000011; // lw    s6,   0(a0)
    assign rom[9'h098] = 32'b00000000010001010010101110000011; // lw    s7,   4(a0)
    assign rom[9'h099] = 32'b00000000100001010010110000000011; // lw    s8,   8(a0)
    assign rom[9'h09a] = 32'b00000000110001010010110010000011; // lw    s9,  12(a0)
    assign rom[9'h09b] = 32'b00000001011010010100100100110011; // xor   s2,  s2,  s6
    assign rom[9'h09c] = 32'b00000001011110011100100110110011; // xor   s3,  s3,  s7
    assign rom[9'h09d] = 32'b00000001100010100100101000110011; // xor   s4,  s4,  s8
    assign rom[9'h09e] = 32'b00000001100110101100101010110011; // xor   s5,  s5,  s9
    assign rom[9'h09f] = 32'b11111111000001010000010100010011; // addi  a0,  a0,  -16
    assign rom[9'h0a0] = 32'b00001111111100000000000110010011; // li    gp,  0xFF
    // aes_dec_block_loop:
    assign rom[9'h0a1] = 32'b00000000001110010111101100110011; // and   s6,   s2,   gp
    assign rom[9'h0a2] = 32'b00000000001110011111101110110011; // and   s7,   s3,   gp
    assign rom[9'h0a3] = 32'b00000000001110100111110000110011; // and   s8,   s4,   gp
    assign rom[9'h0a4] = 32'b00000000001110101111110010110011; // and   s9,   s5,   gp
    assign rom[9'h0a5] = 32'b00000000100000011001110100010011; // slli  s10,  gp,   0x8
    assign rom[9'h0a6] = 32'b00000001101010101111110110110011; // and   s11,  s5,   s10
    assign rom[9'h0a7] = 32'b00000001101110110110101100110011; // or    s6,   s6,   s11
    assign rom[9'h0a8] = 32'b00000001101010010111110110110011; // and   s11,  s2,   s10
    assign rom[9'h0a9] = 32'b00000001101110111110101110110011; // or    s7,   s7,   s11
    assign rom[9'h0aa] = 32'b00000001101010011111110110110011; // and   s11,  s3,   s10
    assign rom[9'h0ab] = 32'b00000001101111000110110000110011; // or    s8,   s8,   s11
    assign rom[9'h0ac] = 32'b00000001101010100111110110110011; // and   s11,  s4,   s10
    assign rom[9'h0ad] = 32'b00000001101111001110110010110011; // or    s9,   s9,   s11
    assign rom[9'h0ae] = 32'b00000000100011010001110100010011; // slli  s10,  s10,  0x8
    assign rom[9'h0af] = 32'b00000001101010100111110110110011; // and   s11,  s4,   s10
    assign rom[9'h0b0] = 32'b00000001101110110110101100110011; // or    s6,   s6,   s11
    assign rom[9'h0b1] = 32'b00000001101010101111110110110011; // and   s11,  s5,   s10
    assign rom[9'h0b2] = 32'b00000001101110111110101110110011; // or    s7,   s7,   s11
    assign rom[9'h0b3] = 32'b00000001101010010111110110110011; // and   s11,  s2,   s10
    assign rom[9'h0b4] = 32'b00000001101111000110110000110011; // or    s8,   s8,   s11
    assign rom[9'h0b5] = 32'b00000001101010011111110110110011; // and   s11,  s3,   s10
    assign rom[9'h0b6] = 32'b00000001101111001110110010110011; // or    s9,   s9,   s11
    assign rom[9'h0b7] = 32'b00000000100011010001110100010011; // slli  s10,  s10,  0x8
    assign rom[9'h0b8] = 32'b00000001101010011111110110110011; // and   s11,  s3,   s10
    assign rom[9'h0b9] = 32'b00000001101110110110101100110011; // or    s6,   s6,   s11
    assign rom[9'h0ba] = 32'b00000001101010100111110110110011; // and   s11,  s4,   s10
    assign rom[9'h0bb] = 32'b00000001101110111110101110110011; // or    s7,   s7,   s11
    assign rom[9'h0bc] = 32'b00000001101010101111110110110011; // and   s11,  s5,   s10
    assign rom[9'h0bd] = 32'b00000001101111000110110000110011; // or    s8,   s8,   s11
    assign rom[9'h0be] = 32'b00000001101010010111110110110011; // and   s11,  s2,   s10
    assign rom[9'h0bf] = 32'b00000001101111001110110010110011; // or    s9,   s9,   s11
    assign rom[9'h0c0] = 32'b00000010000010110001100101111111; // invsubbytes  s2,  s6
    assign rom[9'h0c1] = 32'b00000010000010111001100111111111; // invsubbytes  s3,  s7
    assign rom[9'h0c2] = 32'b00000010000011000001101001111111; // invsubbytes  s4,  s8
    assign rom[9'h0c3] = 32'b00000010000011001001101011111111; // invsubbytes  s5,  s9
    assign rom[9'h0c4] = 32'b00000000000001010010101100000011; // lw   s6,   0(a0)
    assign rom[9'h0c5] = 32'b00000000010001010010101110000011; // lw   s7,   4(a0)
    assign rom[9'h0c6] = 32'b00000000100001010010110000000011; // lw   s8,   8(a0)
    assign rom[9'h0c7] = 32'b00000000110001010010110010000011; // lw   s9,  12(a0)
    assign rom[9'h0c8] = 32'b00000001011010010100100100110011; // xor  s2,  s2,  s6
    assign rom[9'h0c9] = 32'b00000001011110011100100110110011; // xor  s3,  s3,  s7
    assign rom[9'h0ca] = 32'b00000001100010100100101000110011; // xor  s4,  s4,  s8
    assign rom[9'h0cb] = 32'b00000001100110101100101010110011; // xor  s5,  s5,  s9    
    assign rom[9'h0cc] = 32'b00000100000010010001100101111111; // invmixColumns  s2,  s2
    assign rom[9'h0cd] = 32'b00000100000010011001100111111111; // invmixColumns  s3,  s3
    assign rom[9'h0ce] = 32'b00000100000010100001101001111111; // invmixColumns  s4,  s4
    assign rom[9'h0cf] = 32'b00000100000010101001101011111111; // invmixColumns  s5,  s5
    assign rom[9'h0d0] = 32'b11111111000001010000010100010011; // addi  a0,  a0,  -16
    assign rom[9'h0d1] = 32'b11110101000001010001000011100011; // bne a0, a6, aes_dec_block_loop
    // aes_dec_block_finish:
    assign rom[9'h0d2] = 32'b00000000001110010111101100110011; // and   s6,   s2,   gp
    assign rom[9'h0d3] = 32'b00000000001110011111101110110011; // and   s7,   s3,   gp
    assign rom[9'h0d4] = 32'b00000000001110100111110000110011; // and   s8,   s4,   gp
    assign rom[9'h0d5] = 32'b00000000001110101111110010110011; // and   s9,   s5,   gp
    assign rom[9'h0d6] = 32'b00000000100000011001110100010011; // slli  s10,  gp,   0x8
    assign rom[9'h0d7] = 32'b00000001101010101111110110110011; // and   s11,  s5,   s10
    assign rom[9'h0d8] = 32'b00000001101110110110101100110011; // or    s6,   s6,   s11
    assign rom[9'h0d9] = 32'b00000001101010010111110110110011; // and   s11,  s2,   s10
    assign rom[9'h0da] = 32'b00000001101110111110101110110011; // or    s7,   s7,   s11
    assign rom[9'h0db] = 32'b00000001101010011111110110110011; // and   s11,  s3,   s10
    assign rom[9'h0dc] = 32'b00000001101111000110110000110011; // or    s8,   s8,   s11
    assign rom[9'h0dd] = 32'b00000001101010100111110110110011; // and   s11,  s4,   s10
    assign rom[9'h0de] = 32'b00000001101111001110110010110011; // or    s9,   s9,   s11
    assign rom[9'h0df] = 32'b00000000100011010001110100010011; // slli  s10,  s10,  0x8
    assign rom[9'h0e0] = 32'b00000001101010100111110110110011; // and   s11,  s4,   s10
    assign rom[9'h0e1] = 32'b00000001101110110110101100110011; // or    s6,   s6,   s11
    assign rom[9'h0e2] = 32'b00000001101010101111110110110011; // and   s11,  s5,   s10
    assign rom[9'h0e3] = 32'b00000001101110111110101110110011; // or    s7,   s7,   s11
    assign rom[9'h0e4] = 32'b00000001101010010111110110110011; // and   s11,  s2,   s10
    assign rom[9'h0e5] = 32'b00000001101111000110110000110011; // or    s8,   s8,   s11
    assign rom[9'h0e6] = 32'b00000001101010011111110110110011; // and   s11,  s3,   s10
    assign rom[9'h0e7] = 32'b00000001101111001110110010110011; // or    s9,   s9,   s11
    assign rom[9'h0e8] = 32'b00000000100011010001110100010011; // slli  s10,  s10,  0x8
    assign rom[9'h0e9] = 32'b00000001101010011111110110110011; // and   s11,  s3,   s10
    assign rom[9'h0ea] = 32'b00000001101110110110101100110011; // or    s6,   s6,   s11
    assign rom[9'h0eb] = 32'b00000001101010100111110110110011; // and   s11,  s4,   s10
    assign rom[9'h0ec] = 32'b00000001101110111110101110110011; // or    s7,   s7,   s11
    assign rom[9'h0ed] = 32'b00000001101010101111110110110011; // and   s11,  s5,   s10
    assign rom[9'h0ee] = 32'b00000001101111000110110000110011; // or    s8,   s8,   s11
    assign rom[9'h0ef] = 32'b00000001101010010111110110110011; // and   s11,  s2,   s10
    assign rom[9'h0f0] = 32'b00000001101111001110110010110011; // or    s9,   s9,   s11    
    assign rom[9'h0f1] = 32'b00000010000010110001100101111111; // invsubbytes  s2,  s6
    assign rom[9'h0f2] = 32'b00000010000010111001100111111111; // invsubbytes  s3,  s7
    assign rom[9'h0f3] = 32'b00000010000011000001101001111111; // invsubbytes  s4,  s8
    assign rom[9'h0f4] = 32'b00000010000011001001101011111111; // invsubbytes  s5,  s9
    assign rom[9'h0f5] = 32'b00000000000001010010101100000011; // lw   s6,   0(a0)
    assign rom[9'h0f6] = 32'b00000000010001010010101110000011; // lw   s7,   4(a0)
    assign rom[9'h0f7] = 32'b00000000100001010010110000000011; // lw   s8,   8(a0)
    assign rom[9'h0f8] = 32'b00000000110001010010110010000011; // lw   s9,  12(a0)
    assign rom[9'h0f9] = 32'b00000001011010010100100100110011; // xor  s2,  s2,  s6
    assign rom[9'h0fa] = 32'b00000001011110011100100110110011; // xor  s3,  s3,  s7
    assign rom[9'h0fb] = 32'b00000001100010100100101000110011; // xor  s4,  s4,  s8
    assign rom[9'h0fc] = 32'b00000001100110101100101010110011; // xor  s5,  s5,  s9
    assign rom[9'h0fd] = 32'b00000011100000000000100010010011; // la   a7,  output_block
    assign rom[9'h0fe] = 32'b00000001001010001010000000100011; // sw   s2,   0(a7)
    assign rom[9'h0ff] = 32'b00000001001110001010001000100011; // sw   s3,   4(a7)
    assign rom[9'h100] = 32'b00000001010010001010010000100011; // sw   s4,   8(a7)
    assign rom[9'h101] = 32'b00000001010110001010011000100011; // sw   s5,  12(a7)
    assign rom[9'h102] = 32'b00000000000000001000000001100111; // jr   ra
    assign rom[9'h103] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h104] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h105] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h106] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h107] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h108] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h109] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h10a] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h10b] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h10c] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h10d] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h10e] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h10f] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h110] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h111] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h112] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h113] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h114] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h115] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h116] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h117] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h118] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h119] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h11a] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h11b] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h11c] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h11d] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h11e] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h11f] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h120] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h121] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h122] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h123] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h124] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h125] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h126] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h127] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h128] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h129] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h12a] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h12b] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h12c] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h12d] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h12e] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h12f] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h130] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h131] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h132] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h133] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h134] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h135] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h136] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h137] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h138] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h139] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h13a] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h13b] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h13c] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h13d] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h13e] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h13f] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h140] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h141] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h142] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h143] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h144] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h145] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h146] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h147] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h148] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h149] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h14a] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h14b] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h14c] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h14d] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h14e] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h14f] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h150] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h151] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h152] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h153] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h154] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h155] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h156] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h157] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h158] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h159] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h15a] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h15b] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h15c] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h15d] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h15e] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h15f] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h160] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h161] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h162] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h163] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h164] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h165] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h166] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h167] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h168] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h169] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h16a] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h16b] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h16c] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h16d] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h16e] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h16f] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h170] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h171] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h172] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h173] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h174] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h175] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h176] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h177] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h178] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h179] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h17a] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h17b] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h17c] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h17d] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h17e] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h17f] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h180] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h181] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h182] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h183] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h184] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h185] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h186] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h187] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h188] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h189] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h18a] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h18b] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h18c] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h18d] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h18e] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h18f] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h190] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h191] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h192] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h193] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h194] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h195] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h196] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h197] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h198] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h199] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h19a] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h19b] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h19c] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h19d] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h19e] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h19f] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1a0] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1a1] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1a2] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1a3] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1a4] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1a5] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1a6] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1a7] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1a8] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1a9] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1aa] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ab] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ac] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ad] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ae] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1af] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1b0] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1b1] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1b2] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1b3] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1b4] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1b5] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1b6] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1b7] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1b8] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1b9] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ba] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1bb] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1bc] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1bd] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1be] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1bf] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1c0] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1c1] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1c2] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1c3] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1c4] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1c5] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1c6] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1c7] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1c8] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1c9] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ca] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1cb] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1cc] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1cd] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ce] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1cf] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1d0] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1d1] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1d2] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1d3] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1d4] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1d5] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1d6] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1d7] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1d8] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1d9] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1da] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1db] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1dc] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1dd] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1de] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1df] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1e0] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1e1] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1e2] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1e3] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1e4] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1e5] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1e6] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1e7] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1e8] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1e9] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ea] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1eb] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ec] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ed] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ee] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ef] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1f0] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1f1] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1f2] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1f3] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1f4] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1f5] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1f6] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1f7] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1f8] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1f9] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1fa] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1fb] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1fc] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1fd] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1fe] = 32'b00000000000000000000000000000000; // 
    assign rom[9'h1ff] = 32'b00000000000000000000000000000000; // 
    assign inst = rom[a[10:2]];
endmodule